// Code your design here
`include "i2c_master.sv"