`include "simple_if.sv"
`include "tb.sv"