`include "i2c_master.sv"
`include "i2c_slave.sv"