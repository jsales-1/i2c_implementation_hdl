// Code your testbench here
// or browse Examples

`include "i2c_if.sv"
`include "tb.sv"
