// Code your design here
`include "i2c_slave.sv"