`include "assertions.sv"
`include "i2c_tb.sv"